interface xgemac_clk_interface();
    logic clk;

    initial begin
        $display("This is clk interface");
    end
endinterface : xgemac_clk_interface
